// ******************************************************************* //
//                               DEFINE                                //
// ******************************************************************* //

`define DEFAULT_PC   'd0

`define ALU_OP_WIDTH 14

// ******************************************************************* //
//                              LoongArch                              //
// ******************************************************************* //

`define LA64_PC_WIDTH   32
`define LA64_INST_WIDTH 32

`define LA64_ADDR_WIDTH 32
`define LA64_DATA_WIDTH 32

`define LA64_ARF_SEL    5
`define LA64_ARF_NUM    32

